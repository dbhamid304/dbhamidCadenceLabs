* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : OpAmp                                        *
* Netlisted  : Sun Aug 11 22:59:34 2024                     *
* Pegasus Version: 23.20-p013 Tue Jan 9 12:32:47 PST 2024   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n2svt) _nmos_25 ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p2svt) _pmos2v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)
*.DEVTMPLT 2 MP(g45pcap2) _pmoscap2v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369281                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369281 G D_drain_1 B_botTap S_source_0
** N=4 EP=4 FDC=1
M0 D_drain_1 G S_source_0 B_botTap g45n2svt L=7.5e-07 W=6.88e-06 AD=1.032e-12 AS=1.032e-12 PD=1.406e-05 PS=1.406e-05 fw=6.88e-06 sa=1.5e-07 sb=1.5e-07 sca=2.46784 scb=0.000811353 scc=6.29682e-06 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369281

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369282                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369282 G S_source_1 B_botTap D_drain_0
** N=4 EP=4 FDC=1
M0 S_source_1 G D_drain_0 B_botTap g45n2svt L=1.5e-07 W=1.09e-06 AD=1.635e-13 AS=1.635e-13 PD=2.48e-06 PS=2.48e-06 fw=1.09e-06 sa=1.5e-07 sb=1.5e-07 sca=2.69607 scb=5.8866e-05 scc=1.55926e-09 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369282

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmoscap2v_CDNS_723397369283                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmoscap2v_CDNS_723397369283 S_source_0 G D_drain_1 B_tapRight
** N=5 EP=4 FDC=1
M0 D_drain_1 G S_source_0 B_tapRight g45pcap2 L=6.315e-06 W=6.315e-06 AD=9.4725e-13 AS=9.4725e-13 PD=1.293e-05 PS=1.293e-05 $X=0 $Y=0 $dt=2
.ends pmoscap2v_CDNS_723397369283

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_723397369284                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_723397369284 B_topTap G D_drain_1
** N=4 EP=3 FDC=1
M0 D_drain_1 G B_topTap B_topTap g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=9.3e-14 PD=1.33e-06 PS=1.33e-06 fw=4.65e-07 sa=2e-06 sb=1.1e-06 sca=8.22508 scb=0.00662596 scc=0.000256612 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_723397369284

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369285                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369285 D_drain_1 B_botTap 3 4
** N=4 EP=4 FDC=1
M0 D_drain_1 3 4 B_botTap g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=3e-13 PD=3.4e-06 PS=3.4e-06 fw=1.5e-06 sa=2e-06 sb=1.1e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369285

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369286                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369286 G S_source_0 B_botTap 4
** N=4 EP=4 FDC=1
M0 4 G S_source_0 B_botTap g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=3e-13 PD=3.4e-06 PS=3.4e-06 fw=1.5e-06 sa=2e-06 sb=1.1e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369286

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369287                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369287 D_drain_1 G S_source_0 B_botTap
** N=4 EP=4 FDC=1
M0 D_drain_1 G S_source_0 B_botTap g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=2.25e-13 PD=3.4e-06 PS=3.3e-06 fw=1.5e-06 sa=1.5e-07 sb=2e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369287

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_723397369288                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_723397369288 B_topTap S_source_0 G
** N=4 EP=3 FDC=1
M0 G G S_source_0 B_topTap g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=6.975e-14 PD=1.33e-06 PS=1.23e-06 fw=4.65e-07 sa=1.5e-07 sb=2e-06 sca=9.90286 scb=0.00793993 scc=0.000268631 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_723397369288

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369289                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369289 S_source_0 B_botTap 3 4
** N=4 EP=4 FDC=1
M0 4 3 S_source_0 B_botTap g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=2.25e-13 PD=3.4e-06 PS=3.3e-06 fw=1.5e-06 sa=1.5e-07 sb=2e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369289

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_7233973692810                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_7233973692810 B_topTap S_source_0 G D_drain_1
** N=5 EP=4 FDC=1
M0 D_drain_1 G S_source_0 B_topTap g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=6.975e-14 PD=1.33e-06 PS=1.23e-06 fw=4.65e-07 sa=1.5e-07 sb=2e-06 sca=9.90286 scb=0.00793993 scc=0.000268631 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_7233973692810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_7233973692811                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_7233973692811 B_topTap S_source_0 G 4
** N=5 EP=4 FDC=1
M0 4 G S_source_0 B_topTap g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=9.3e-14 PD=1.33e-06 PS=1.33e-06 fw=4.65e-07 sa=2e-06 sb=1.1e-06 sca=8.22508 scb=0.00662596 scc=0.000256612 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_7233973692811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_7233973692812                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_7233973692812 D_drain_0 B_botTap G S_source_1
** N=4 EP=4 FDC=1
M0 S_source_1 G D_drain_0 B_botTap g45n2svt L=7.5e-07 W=1.09e-06 AD=1.635e-13 AS=1.635e-13 PD=2.48e-06 PS=2.48e-06 fw=1.09e-06 sa=1.5e-07 sb=1.5e-07 sca=2.09979 scb=2.24679e-05 scc=4.87113e-10 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_7233973692812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OpAmp                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OpAmp IBIAS INN INP OUT VDD VSS
** N=9 EP=6 FDC=13
X53 IBIAS VSS VSS OUT nmos2v_CDNS_723397369281 $T=20520 18100 0 180 $X=18360 $Y=3980
X54 IBIAS VSS VSS 9 nmos2v_CDNS_723397369282 $T=16430 2540 1 0 $X=15770 $Y=0
X55 OUT 2 OUT OUT pmoscap2v_CDNS_723397369283 $T=3840 21800 1 0 $X=3060 $Y=8690
X56 VDD 8 8 pmos2v_CDNS_723397369284 $T=10110 7010 0 180 $X=7870 $Y=4640
X57 2 VSS INP 9 nmos2v_CDNS_723397369285 $T=10110 3360 0 180 $X=7990 $Y=0
X58 INN 9 VSS 8 nmos2v_CDNS_723397369286 $T=10510 3360 1 0 $X=9890 $Y=0
X59 8 INN 9 VSS nmos2v_CDNS_723397369287 $T=13910 3360 0 180 $X=11790 $Y=0
X60 VDD VDD 8 pmos2v_CDNS_723397369288 $T=6710 7010 1 0 $X=5930 $Y=4640
X61 9 VSS INP 2 nmos2v_CDNS_723397369289 $T=6710 3360 1 0 $X=6050 $Y=0
X62 VDD VDD 8 2 pmos2v_CDNS_7233973692810 $T=13910 7010 0 180 $X=11670 $Y=4640
X63 VDD VDD 8 2 pmos2v_CDNS_7233973692811 $T=10510 7010 1 0 $X=9770 $Y=4640
X64 VSS VSS IBIAS IBIAS nmos2v_CDNS_7233973692812 $T=19020 2540 1 0 $X=18360 $Y=0
M0 OUT 2 VDD VDD g45p2svt L=1.5e-07 W=1e-05 AD=1.5e-12 AS=1.5e-12 PD=2.03e-05 PS=2.03e-05 fw=1e-05 sa=1.5e-07 sb=1.5e-07 sca=10.0331 scb=0.00968513 scc=0.0001241 $X=780 $Y=1560 $dt=1
.ends OpAmp
