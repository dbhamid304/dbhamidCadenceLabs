* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : OpAmp                                        *
* Netlisted  : Sun Aug 11 22:59:34 2024                     *
* Pegasus Version: 23.20-p013 Tue Jan 9 12:32:47 PST 2024   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n2svt) _nmos_25 ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p2svt) _pmos2v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)
*.DEVTMPLT 2 MP(g45pcap2) _pmoscap2v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_723397369280                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_723397369280 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_723397369280

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_723397369282                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_723397369282 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_723397369282

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_723397369283                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_723397369283 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_723397369283

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_723397369284                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_723397369284 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_723397369284

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_723397369285                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_723397369285 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_723397369285

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_723397369286                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_723397369286 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_723397369286

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_723397369287                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_723397369287 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_723397369287

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_723397369289                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_723397369289 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_723397369289

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7233973692810                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7233973692810 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7233973692810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7233973692811                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7233973692811 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7233973692811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7233973692815                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7233973692815 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7233973692815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369281                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369281 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 4 3 g45n2svt L=7.5e-07 W=6.88e-06 AD=1.032e-12 AS=1.032e-12 PD=1.406e-05 PS=1.406e-05 fw=6.88e-06 sa=1.5e-07 sb=1.5e-07 sca=2.46784 scb=0.000811353 scc=6.29682e-06 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369281

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369282                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369282 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 4 3 g45n2svt L=1.5e-07 W=1.09e-06 AD=1.635e-13 AS=1.635e-13 PD=2.48e-06 PS=2.48e-06 fw=1.09e-06 sa=1.5e-07 sb=1.5e-07 sca=2.69607 scb=5.8866e-05 scc=1.55926e-09 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369282

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmoscap2v_CDNS_723397369283                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmoscap2v_CDNS_723397369283 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 4 g45pcap2 L=6.315e-06 W=6.315e-06 AD=9.4725e-13 AS=9.4725e-13 PD=1.293e-05 PS=1.293e-05 $X=0 $Y=0 $dt=2
.ends pmoscap2v_CDNS_723397369283

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_723397369284                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_723397369284 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 1 g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=9.3e-14 PD=1.33e-06 PS=1.33e-06 fw=4.65e-07 sa=2e-06 sb=1.1e-06 sca=8.22508 scb=0.00662596 scc=0.000256612 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_723397369284

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369285                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369285 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 3 4 2 g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=3e-13 PD=3.4e-06 PS=3.4e-06 fw=1.5e-06 sa=2e-06 sb=1.1e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369285

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369286                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369286 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 1 2 3 g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=3e-13 PD=3.4e-06 PS=3.4e-06 fw=1.5e-06 sa=2e-06 sb=1.1e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369286

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369287                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369287 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=2.25e-13 PD=3.4e-06 PS=3.3e-06 fw=1.5e-06 sa=1.5e-07 sb=2e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369287

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_723397369288                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_723397369288 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 3 2 1 g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=6.975e-14 PD=1.33e-06 PS=1.23e-06 fw=4.65e-07 sa=1.5e-07 sb=2e-06 sca=9.90286 scb=0.00793993 scc=0.000268631 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_723397369288

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_723397369289                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_723397369289 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n2svt L=7.5e-07 W=1.5e-06 AD=3e-13 AS=2.25e-13 PD=3.4e-06 PS=3.3e-06 fw=1.5e-06 sa=1.5e-07 sb=2e-06 sca=2.273 scb=9.86043e-05 scc=6.38585e-08 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_723397369289

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_7233973692810                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_7233973692810 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 4 3 2 1 g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=6.975e-14 PD=1.33e-06 PS=1.23e-06 fw=4.65e-07 sa=1.5e-07 sb=2e-06 sca=9.90286 scb=0.00793993 scc=0.000268631 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_7233973692810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos2v_CDNS_7233973692811                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos2v_CDNS_7233973692811 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 4 3 2 1 g45p2svt L=7.5e-07 W=4.65e-07 AD=9.3e-14 AS=9.3e-14 PD=1.33e-06 PS=1.33e-06 fw=4.65e-07 sa=2e-06 sb=1.1e-06 sca=8.22508 scb=0.00662596 scc=0.000256612 $X=0 $Y=0 $dt=1
.ends pmos2v_CDNS_7233973692811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos2v_CDNS_7233973692812                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos2v_CDNS_7233973692812 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n2svt L=7.5e-07 W=1.09e-06 AD=1.635e-13 AS=1.635e-13 PD=2.48e-06 PS=2.48e-06 fw=1.09e-06 sa=1.5e-07 sb=1.5e-07 sca=2.09979 scb=2.24679e-05 scc=4.87113e-10 $X=0 $Y=0 $dt=0
.ends nmos2v_CDNS_7233973692812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OpAmp                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OpAmp 6 4 3 7 1 5
** N=9 EP=6 FDC=13
X0 1 M2_M1_CDNS_723397369280 $T=950 11080 0 0 $X=820 $Y=10950
X1 1 M2_M1_CDNS_723397369280 $T=2340 5670 0 0 $X=2210 $Y=5540
X2 2 M2_M1_CDNS_723397369280 $T=5750 1360 0 0 $X=5620 $Y=1230
X3 3 M2_M1_CDNS_723397369280 $T=6450 3800 0 0 $X=6320 $Y=3670
X4 1 M2_M1_CDNS_723397369280 $T=10310 5240 0 0 $X=10180 $Y=5110
X5 4 M2_M1_CDNS_723397369280 $T=11210 3560 0 0 $X=11080 $Y=3430
X6 1 M2_M1_CDNS_723397369280 $T=14090 5240 0 0 $X=13960 $Y=5110
X7 5 M2_M1_CDNS_723397369280 $T=16910 3380 0 0 $X=16780 $Y=3250
X8 5 M2_M1_CDNS_723397369280 $T=18840 3380 0 0 $X=18710 $Y=3250
X9 5 M2_M1_CDNS_723397369280 $T=18840 18940 0 0 $X=18710 $Y=18810
X10 6 M2_M1_CDNS_723397369280 $T=19890 2740 0 0 $X=19760 $Y=2610
X11 6 M2_M1_CDNS_723397369280 $T=19890 4140 0 0 $X=19760 $Y=4010
X12 7 M3_M2_CDNS_723397369282 $T=16650 18470 0 0 $X=16520 $Y=18220
X13 7 M3_M2_CDNS_723397369282 $T=17610 18470 0 0 $X=17480 $Y=18220
X14 4 M3_M2_CDNS_723397369283 $T=160 4630 0 0 $X=30 $Y=4500
X15 6 M3_M2_CDNS_723397369283 $T=160 8270 0 0 $X=30 $Y=8140
X16 2 M3_M2_CDNS_723397369283 $T=8410 3740 0 0 $X=8280 $Y=3610
X17 8 M3_M2_CDNS_723397369283 $T=8410 5700 0 0 $X=8280 $Y=5570
X18 4 M3_M2_CDNS_723397369283 $T=11210 4630 0 0 $X=11080 $Y=4500
X19 8 M3_M2_CDNS_723397369283 $T=12210 5700 0 0 $X=12080 $Y=5570
X20 7 M3_M2_CDNS_723397369283 $T=21020 18470 0 0 $X=20890 $Y=18340
X21 1 M2_M1_CDNS_723397369284 $T=6530 5240 0 0 $X=6450 $Y=5110
X22 1 M2_M1_CDNS_723397369284 $T=6530 6545 0 0 $X=6450 $Y=6415
X23 2 M2_M1_CDNS_723397369284 $T=8410 2580 0 0 $X=8330 $Y=2450
X24 8 M2_M1_CDNS_723397369284 $T=8410 6080 0 0 $X=8330 $Y=5950
X25 1 M2_M1_CDNS_723397369284 $T=10310 6410 0 0 $X=10230 $Y=6280
X26 8 M2_M1_CDNS_723397369284 $T=12210 2820 0 0 $X=12130 $Y=2690
X27 1 M2_M1_CDNS_723397369284 $T=14090 6390 0 0 $X=14010 $Y=6260
X28 5 M2_M1_CDNS_723397369284 $T=16910 1590 0 0 $X=16830 $Y=1460
X29 5 M2_M1_CDNS_723397369284 $T=18840 1450 0 0 $X=18760 $Y=1320
X30 5 M2_M1_CDNS_723397369284 $T=18840 11220 0 0 $X=18760 $Y=11090
X31 2 M2_M1_CDNS_723397369285 $T=12210 6545 0 0 $X=12130 $Y=6295
X32 7 M2_M1_CDNS_723397369285 $T=16650 18470 0 0 $X=16570 $Y=18220
X33 7 M2_M1_CDNS_723397369285 $T=17610 18470 0 0 $X=17530 $Y=18220
X34 2 M2_M1_CDNS_723397369286 $T=12210 8970 0 0 $X=11960 $Y=8890
X35 6 M2_M1_CDNS_723397369286 $T=19340 2740 0 0 $X=19090 $Y=2660
X36 8 M3_M2_CDNS_723397369287 $T=7460 5700 0 0 $X=7210 $Y=5620
X37 8 M3_M2_CDNS_723397369287 $T=9420 5700 0 0 $X=9170 $Y=5620
X38 8 M3_M2_CDNS_723397369287 $T=11390 5700 0 0 $X=11140 $Y=5620
X39 8 M3_M2_CDNS_723397369287 $T=13120 5700 0 0 $X=12870 $Y=5620
X40 6 M3_M2_CDNS_723397369287 $T=19340 2740 0 0 $X=19090 $Y=2660
X41 7 M3_M2_CDNS_723397369287 $T=20700 18470 0 0 $X=20450 $Y=18390
X42 2 M4_M3_CDNS_723397369289 $T=12210 3740 0 0 $X=12080 $Y=3610
X43 6 M4_M3_CDNS_723397369289 $T=16580 8270 0 0 $X=16450 $Y=8140
X44 2 M3_M2_CDNS_7233973692810 $T=12210 6545 0 0 $X=12130 $Y=6295
X45 6 M3_M2_CDNS_7233973692810 $T=16580 2740 0 0 $X=16500 $Y=2490
X46 2 M4_M3_CDNS_7233973692811 $T=12210 6545 0 0 $X=12130 $Y=6295
X47 6 M4_M3_CDNS_7233973692811 $T=16580 2740 0 0 $X=16500 $Y=2490
X48 8 M2_M1_CDNS_7233973692815 $T=7460 5700 0 0 $X=7210 $Y=5570
X49 8 M2_M1_CDNS_7233973692815 $T=9420 5700 0 0 $X=9170 $Y=5570
X50 8 M2_M1_CDNS_7233973692815 $T=11390 5700 0 0 $X=11140 $Y=5570
X51 8 M2_M1_CDNS_7233973692815 $T=13120 5700 0 0 $X=12870 $Y=5570
X52 7 M2_M1_CDNS_7233973692815 $T=20700 18470 0 0 $X=20450 $Y=18340
X53 6 5 5 7 nmos2v_CDNS_723397369281 $T=20520 18100 0 180 $X=18360 $Y=3980
X54 6 5 5 9 nmos2v_CDNS_723397369282 $T=16430 2540 1 0 $X=15770 $Y=0
X55 7 2 7 7 5 pmoscap2v_CDNS_723397369283 $T=3840 21800 1 0 $X=3060 $Y=8690
X56 1 8 8 5 pmos2v_CDNS_723397369284 $T=10110 7010 0 180 $X=7870 $Y=4640
X57 2 5 3 9 nmos2v_CDNS_723397369285 $T=10110 3360 0 180 $X=7990 $Y=0
X58 4 9 5 8 nmos2v_CDNS_723397369286 $T=10510 3360 1 0 $X=9890 $Y=0
X59 8 4 9 5 nmos2v_CDNS_723397369287 $T=13910 3360 0 180 $X=11790 $Y=0
X60 1 1 8 5 pmos2v_CDNS_723397369288 $T=6710 7010 1 0 $X=5930 $Y=4640
X61 9 5 3 2 nmos2v_CDNS_723397369289 $T=6710 3360 1 0 $X=6050 $Y=0
X62 1 1 8 2 5 pmos2v_CDNS_7233973692810 $T=13910 7010 0 180 $X=11670 $Y=4640
X63 1 1 8 2 5 pmos2v_CDNS_7233973692811 $T=10510 7010 1 0 $X=9770 $Y=4640
X64 5 5 6 6 nmos2v_CDNS_7233973692812 $T=19020 2540 1 0 $X=18360 $Y=0
M0 7 2 1 1 g45p2svt L=1.5e-07 W=1e-05 AD=1.5e-12 AS=1.5e-12 PD=2.03e-05 PS=2.03e-05 fw=1e-05 sa=1.5e-07 sb=1.5e-07 sca=10.0331 scb=0.00968513 scc=0.0001241 $X=780 $Y=1560 $dt=1
.ends OpAmp
